architecture btnMode_a of btnMode_e is

  type mode_st is (mode2_st, mode3_st, mode4_st, mode5_st);

begin


